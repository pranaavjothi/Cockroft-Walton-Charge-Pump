* C:\Users\prana\eSim-Workspace\cockroft_walton_charge_pump\cockroft_walton_charge_pump.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/04/22 12:05:29

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  GND GND Net-_C1-Pad1_ GND eSim_MOS_N		
M2  Net-_C1-Pad1_ Net-_C1-Pad1_ Net-_C2-Pad1_ GND eSim_MOS_N		
M3  Net-_C2-Pad1_ Net-_C2-Pad1_ Net-_C3-Pad1_ GND eSim_MOS_N		
M4  Net-_C3-Pad1_ Net-_C3-Pad1_ out GND eSim_MOS_N		
C1  Net-_C1-Pad1_ in 1u		
C2  Net-_C2-Pad1_ GND 1u		
C3  Net-_C3-Pad1_ Net-_C1-Pad1_ 1u		
C4  out Net-_C2-Pad1_ 1u		
U1  in plot_v1		
U2  out plot_v1		
v1  in GND sine		

.end
